-------------------------------------------------
--  File:          haC64.vhd
--
--  Entity:        haC64
--  Architecture:  Structural
--  Author:        Seth Gower and Paul Kelly
--  Created:       02/16/19
--  Modified:      
--  VHDL'93
--  Description:   The following is the entity and
--                 architectural description of a
--                 Commodore 64 for BrickHack V at
--                 RIT
-------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity haC64 is
    port(
        clk     : in    std_logic
    );
end entity haC64;
architecture Structural of haC64 is
begin
end Structural;
