-------------------------------------------------
--  File:          name.vhd
--
--  Entity:        entity
--  Architecture:  arch
--  Author:        Seth Gower and Paul Kelly
--  Created:       02/16/19
--  Modified:      
--  VHDL'93
--  Description:   
-------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity ent is
    port(
        clk     : in    std_logic
    );
end entity ent;
architecture arch of ent is
begin
end arch;
